-- Copyright (C) 2012 Carla Sauvanaud
-- Copyright (C) 2012, 2016  Benoît Morgan
--
-- This file is part of dumb8.
--
-- dumb8 is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- dumb8 is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with dumb8.  If not, see <http://www.gnu.org/licenses/>.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity op_to_rw_memoire_donnees is
    Port ( Op : in  STD_LOGIC_VECTOR (7 downto 0);
           RW : out  STD_LOGIC);
end op_to_rw_memoire_donnees;

architecture Behavioral of op_to_rw_memoire_donnees is

begin

with Op select
	RW <= '0' when x"08",
			  '1' when others;

end Behavioral;

