// OP codes
parameter OP_ADD = 8'h01;
parameter OP_SOU = 8'h02;
parameter OP_SHL = 8'h03;
parameter OP_SHR = 8'h04;
parameter OP_COP = 8'h05;
parameter OP_AFC = 8'h06;
parameter OP_LOD = 8'h07;
parameter OP_STR = 8'h08;
parameter OP_JMP = 8'h09;
parameter OP_JMZ = 8'h0A;
