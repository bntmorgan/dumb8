/*
Copyright (C) 2012 Carla Sauvanaud
Copyright (C) 2012, 2016  Benoît Morgan

This file is part of dumb8.

dumb8 is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

dumb8 is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with dumb8.  If not, see <http://www.gnu.org/licenses/>.
*/

// OP codes
parameter OP_ADD = 8'h01;
parameter OP_SOU = 8'h02;
parameter OP_SHL = 8'h03;
parameter OP_SHR = 8'h04;
parameter OP_COP = 8'h05;
parameter OP_AFC = 8'h06;
parameter OP_LOD = 8'h07;
parameter OP_STR = 8'h08;
parameter OP_JMP = 8'h09;
parameter OP_JMZ = 8'h0a;
parameter OP_VWR = 8'h0b;
